library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package serpent_pkg is
end package serpent_pkg;

package body serpent_pkg is
end package body;