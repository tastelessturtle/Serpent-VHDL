library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity serpent is
end entity serpent;

architecture rtl of serpent is
begin
end architecture rtl;